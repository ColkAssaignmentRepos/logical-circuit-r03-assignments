module m_adder(input [3:0] in1, input [3:0] in2, output [7:0] result);
	assign result = in1 + in2;
endmodule
